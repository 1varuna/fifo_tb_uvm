// Package cannot include Interface file!!
package fifo_rtl_pkg;
	
	`include "fifo.sv"	

endpackage
