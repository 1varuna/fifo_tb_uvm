`define DEF_FIFO_WIDTH 32
`define DEF_FIFO_DEPTH 2**5
